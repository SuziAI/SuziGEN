BZh91AY&SY�|�M '߀Py���������`�m�3�    t t7m���     �#i43H�1@2b�d2@jz
�  @��� 9�#� �&���0F&�����1 ѧ�  i��  $�4��SdG���4�SL�cBzA"h����ɣF�4@Y���QD�F����	
���$(���	!GT5��)RI?W�"�I<fUʈgӼrG���l� o����#�(�8*0��#��@$i����f..ۥV��&V�	mLKr��`�2*0��`ك.��	pqq���`@���fƒڡ ��}y�9	�E�?P��-�|��0ߺ��Cj��8HX(`K�	�HA��:36�ܠ��V�5TV�{�wB�j�ɰ�\T-�9.^(�'L
�R/(�iTә����6uvDM9e�as':D8��=�{A��4NT��`58Y���BYf(�Kɺ7jn�m[Z�H�������Dz�&��+st���(q���KC��Jڕ� �N���D�Y�J��������0�z�N��Ƴ��ӏ%$��d�,��S0�fApbKP�(�75oq8,;UF���Y�2�� M�(qÑ��Z�� ��k�U�nJ+ĸ'h���~���_.�n��n3!pѱ�>�`a����KAF�G7aae����`<��A�و�ޗ9�)���!���²�р��^�N��a��a���1`�P�E�c����R9iASw���j�E@�BBp�}��������9meψ����dssp,c�Q&�tA%2�"�:�w�(L�[e�A�QN���T���X�\V$6�V����i�o��!��s�<;���_>�����iB��|��!���)5|����lWl+����)4H�ᮆ��	Y�F�E��I/���#"��
,sZq���D���&f-�r�	��@���´��.�rQj6��5�Y#���"=4�V[���OvC�PC��Ԡ:[���!#Й�>�`<1�����AP䉀�D��B%�5��h�G��Bz����n�z�Uӌ�TD���P0a�4�5��>�ܸ	kB�0d�8P{ADI�	��B�e������Nh�W�48�m�38܅4p4{d�"%�q+�����e
D�l��[ "��J� Nwk ��~��>s@�Ϡ�	0`�C�:��ڱ}0����C�$9&����$,��I� :����2L49�!&l([�,�1B�qi��GN�5򗔪�nl�����0�6I$ʻ���G�>�JKs|QSQrG�S.��Z�Ä�tJ�`]��|���)t�g0����vl,F�a���<9VI�eyT��6�f3�|fZ�i`3aA��t��Á���O�E{xYӴO+;���.&������u��?'6ci�5+GǖP|�Ja4-TI�a<���RZa���4\#b���aY���-Gt��-�Q�~rJ���կ�����g~*��ń�{"�MkAD@X]Յ�J�ʬ�Uh�.B9FT=�|<���#���\[�cl�j'G?-������t-�3m�i���Oy����$a��Y;}�8�7Xt�"MVA`Ý����
�7����m�{V����:��=*��Hf�wڠ�{h�E�e���s��:��f�����N;d��EU���rI$}�t4B���PB�ݜ<p��d��)�PL	�N�X�B��.B6Җ���6�ڰ���Eh��#m����nr�w�����q�G�h��:�����bn�z��.�R��[%���0�%��9~�,m�/�������A���|�0X1�k��a��5���qp�u��}��z�xxɘ\���g-�W�ߡhDF��UUU�	D}�q�r'Ҹ�G� ��0��8|.
G�BE�Oh�8PQ�ʜH��J�i����
��]XE+KE#CE+IEKh�+!�����--U
 ���`SI�-0�&&-�@�cl �YȔ�"H��%����F���� �i*�I� ƃ���@u�Ų�G+���u��	�Jg�q�����$�H�ؘ�#V�v��L�yŵ���
� 
`�k�NIr>�M�TQva� @�^o����'���M-e
kY��q�X��}	�����Ì��.��`�⻏f�������| ��CR�E@��K%	�S�j}$0�yv�!�&"{V%�)���e���l�R���P3���?�y!�b%'DD޴���C\pX0��1_��%%'�2����ҕ{�|`+��q4�Cn8%�aE�#���Lz��[�얅��"%��Q�*�@��0�$ 0 @W+\�T���e��!�S�_���z.iV!���;��{M��(�"��Z"�*��ܮ>��:9X���3|B؛�4A�[�}q&���=�rW �Z&��1������9��P):��"�e`�#�z�����/�=?C�:4�d��`w��zc�����N ��} |��H����|7V�����sټzD7l�p�D�)Z����kg�[M2�P��b��QB��+����4�,�2���eBsX���ȱ�.�t
m ���v�\rB�BY߀G@/�k�*�	�ng�S�1S3!�S� ��%��"+�Jh9�T�MKw#zض�8}�-��Lᘞ��B�� 3����:8-�P>�Oo�]���Jo�Q\)�Q�߬=�grzN5��A�n�P�.r��-�u$=BpH#�R{���N-�h�4DT
]H����>��E@���C���+��xV��z�V����7߈8����c�(�b���I�w6+���'1ѠvkV��;3�%��v.���ji��.���DLw��׎%J((�Iƛ��������N���\�E<4tH K�ݙ`��2�9Ev�G�7����"��b��{��"�ANPW�q�o�k3��n����8�?�*��*^9�������*�;R	o�z���.�p�!H���